

module activation_unit(
	input clk,
	input rstn,	
	input type [2:0]
);

	// Quantize into activation type
	// ReLU, tanh, e 

endmodule

