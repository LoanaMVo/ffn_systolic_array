// RELU
//McMaster Universiry, 4OJ4 Individual Research Course
// Author: Loana
// Date: Febuary 2024
module relu #(
    parameter DATA_WIDTH = 8
)(
    input logic signed  [DATA_WIDTH-1:0] z_i,
    output logic signed [DATA_WIDTH-1:0] y_o
);
always_comb: begin
    if(|z_i[DATA_WIDTH-1]) y_o = '0; // check MSB for negative
    else begin
        case(z_i):
            8'd0   : y_o = 8'b00000000;
            8'd1   : y_o = 8'b00000001;
            8'd2   : y_o = 8'b00000010;
            8'd3   : y_o = 8'b00000011;
            8'd4   : y_o = 8'b00000100;
            8'd5   : y_o = 8'b00000101;
            8'd6   : y_o = 8'b00000110;
            8'd7   : y_o = 8'b00000111;
            8'd8   : y_o = 8'b00001000;
            8'd9   : y_o = 8'b00001001;
            8'd10  : y_o = 8'b00001010;
            8'd11  : y_o = 8'b00001011;
            8'd12  : y_o = 8'b00001100;
            8'd13  : y_o = 8'b00001101;
            8'd14  : y_o = 8'b00001110;
            8'd15  : y_o = 8'b00001111;
            8'd16  : y_o = 8'b00010000;
            8'd17  : y_o = 8'b00010001;
            8'd18  : y_o = 8'b00010010;
            8'd19  : y_o = 8'b00010011;
            8'd20  : y_o = 8'b00010100;
            8'd21  : y_o = 8'b00010101;
            8'd22  : y_o = 8'b00010110;
            8'd23  : y_o = 8'b00010111;
            8'd24  : y_o = 8'b00011000;
            8'd25  : y_o = 8'b00011001;
            8'd26  : y_o = 8'b00011010;
            8'd27  : y_o = 8'b00011011;
            8'd28  : y_o = 8'b00011100;
            8'd29  : y_o = 8'b00011101;
            8'd30  : y_o = 8'b00011110;
            8'd31  : y_o = 8'b00011111;
            8'd32  : y_o = 8'b00100000;
            8'd33  : y_o = 8'b00100001;
            8'd34  : y_o = 8'b00100010;
            8'd35  : y_o = 8'b00100011;
            8'd36  : y_o = 8'b00100100;
            8'd37  : y_o = 8'b00100101;
            8'd38  : y_o = 8'b00100110;
            8'd39  : y_o = 8'b00100111;
            8'd40  : y_o = 8'b00101000;
            8'd41  : y_o = 8'b00101001;
            8'd42  : y_o = 8'b00101010;
            8'd43  : y_o = 8'b00101011;
            8'd44  : y_o = 8'b00101100;
            8'd45  : y_o = 8'b00101101;
            8'd46  : y_o = 8'b00101110;
            8'd47  : y_o = 8'b00101111;
            8'd48  : y_o = 8'b00110000;
            8'd49  : y_o = 8'b00110001;
            8'd50  : y_o = 8'b00110010;
            8'd51  : y_o = 8'b00110011;
            8'd52  : y_o = 8'b00110100;
            8'd53  : y_o = 8'b00110101;
            8'd54  : y_o = 8'b00110110;
            8'd55  : y_o = 8'b00110111;
            8'd56  : y_o = 8'b00111000;
            8'd57  : y_o = 8'b00111001;
            8'd58  : y_o = 8'b00111010;
            8'd59  : y_o = 8'b00111011;
            8'd60  : y_o = 8'b00111100;
            8'd61  : y_o = 8'b00111101;
            8'd62  : y_o = 8'b00111110;
            8'd63  : y_o = 8'b00111111;
            8'd64  : y_o = 8'b01000000;
            8'd65  : y_o = 8'b01000001;
            8'd66  : y_o = 8'b01000010;
            8'd67  : y_o = 8'b01000011;
            8'd68  : y_o = 8'b01000100;
            8'd69  : y_o = 8'b01000101;
            8'd70  : y_o = 8'b01000110;
            8'd71  : y_o = 8'b01000111;
            8'd72  : y_o = 8'b01001000;
            8'd73  : y_o = 8'b01001001;
            8'd74  : y_o = 8'b01001010;
            8'd75  : y_o = 8'b01001011;
            8'd76  : y_o = 8'b01001100;
            8'd77  : y_o = 8'b01001101;
            8'd78  : y_o = 8'b01001110;
            8'd79  : y_o = 8'b01001111;
            8'd80  : y_o = 8'b01010000;
            8'd81  : y_o = 8'b01010001;
            8'd82  : y_o = 8'b01010010;
            8'd83  : y_o = 8'b01010011;
            8'd84  : y_o = 8'b01010100;
            8'd85  : y_o = 8'b01010101;
            8'd86  : y_o = 8'b01010110;
            8'd87  : y_o = 8'b01010111;
            8'd88  : y_o = 8'b01011000;
            8'd89  : y_o = 8'b01011001;
            8'd90  : y_o = 8'b01011010;
            8'd91  : y_o = 8'b01011011;
            8'd92  : y_o = 8'b01011100;
            8'd93  : y_o = 8'b01011101;
            8'd94  : y_o = 8'b01011110;
            8'd95  : y_o = 8'b01011111;
            8'd96  : y_o = 8'b01100000;
            8'd97  : y_o = 8'b01100001;
            8'd98  : y_o = 8'b01100010;
            8'd99  : y_o = 8'b01100011;
            8'd100 : y_o = 8'b01100100;
            8'd101 : y_o = 8'b01100101;
            8'd102 : y_o = 8'b01100110;
            8'd103 : y_o = 8'b01100111;
            8'd104 : y_o = 8'b01101000;
            8'd105 : y_o = 8'b01101001;
            8'd106 : y_o = 8'b01101010;
            8'd107 : y_o = 8'b01101011;
            8'd108 : y_o = 8'b01101100;
            8'd109 : y_o = 8'b01101101;
            8'd110 : y_o = 8'b01101110;
            8'd111 : y_o = 8'b01101111;
            8'd112 : y_o = 8'b01110000;
            8'd113 : y_o = 8'b01110001;
            8'd114 : y_o = 8'b01110010;
            8'd115 : y_o = 8'b01110011;
            8'd116 : y_o = 8'b01110100;
            8'd117 : y_o = 8'b01110101;
            8'd118 : y_o = 8'b01110110;
            8'd119 : y_o = 8'b01110111;
            8'd120 : y_o = 8'b01111000;
            8'd121 : y_o = 8'b01111001;
            8'd122 : y_o = 8'b01111010;
            8'd123 : y_o = 8'b01111011;
            8'd124 : y_o = 8'b01111100;
            8'd125 : y_o = 8'b01111101;
            8'd126 : y_o = 8'b01111110;
            8'd127 : y_o = 8'b01111111;
        endcase
    end
end
endmodule //relu